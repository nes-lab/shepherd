** Profile: "SCHEMATIC1-simIlate"  [ C:\Users\ingmo\Documents\GitHub\shepherd_v2_planning\PCBs\shepherd_recorder_opDrain-PSpiceFiles\SCHEMATIC1\simIlate.sim ]

** Creating circuit file "simIlate.cir"
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries:
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib"
.lib "nom.lib"

*Analysis directives:
.TRAN  0 0.01 0
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*))
.INC "..\SCHEMATIC1.net"


.END
